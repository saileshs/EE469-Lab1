library verilog;
use verilog.vl_types.all;
entity nor_testbench is
end nor_testbench;
