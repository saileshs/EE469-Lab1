library verilog;
use verilog.vl_types.all;
entity cpu_testbench is
end cpu_testbench;
