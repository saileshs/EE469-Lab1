library verilog;
use verilog.vl_types.all;
entity SE_testbench is
end SE_testbench;
