library verilog;
use verilog.vl_types.all;
entity controlUnit_testbench is
end controlUnit_testbench;
