library verilog;
use verilog.vl_types.all;
entity decoder_testbench is
end decoder_testbench;
