library verilog;
use verilog.vl_types.all;
entity mux_testbench is
end mux_testbench;
